module filler( b,a);
  input  [36:1] a;
  output reg [36:1] b;
  wire [6:1] sum;
  assign sum=a[4:1]+ a[8:5]+ a[12:9]+ a[16:13]+ a[20:17]+ a[24:21]+ a[28:25]+a[32:29]+ a[36:33] ;
  always @(a)begin
  case (  { !a[36:33],!a[32:29],!a[28:25],!a[24:21],!a[20:17],!a[16:13],!a[12:9],!a[8:5],!a[4:1]}  )
    9'd1: begin
             b[4:1]= 6'd45 - sum;
             b[36:5]<=a[36:5];
            
           end
    9'd2: begin
      b[8:5]= 6'd45 - sum;
      b[36:9]<=a[36:9];
      b[4:1]<=a[4:1];
    end
     9'd4: begin
       b[12:9]= 6'd45 - sum;
       b[36:13]<=a[36:13];
       b[8:1]<=a[8:1];
    end
     9'd8: begin
       b[16:13]= 6'd45 - sum;
       b[36:17]<=a[36:17];
       b[12:1]<=a[12:1];
    end
     9'd16 : begin
       b[20:17]= 6'd45 - sum;
       b[36:21]<=a[36:21];
       b[16:1]<=a[16:1];
    end
    
     9'b000100000 : begin
       b[24:21]= 6'd45 - sum;
       b[36:25]<=a[36:25];
       b[20:1]<=a[20:1];
    end
    9'b001000000 : begin
      b[28:25]= 6'd45 - sum;
      b[36:29]<=a[36:29];
      b[24:1]<=a[24:1];
    end
    9'b010000000 : begin
      b[32:29]= 6'd45 - sum;
      b[36:33]<=a[36:33];
      b[28:1]<=a[28:1];
    end
     9'b100000000 : begin
       b[36:33]= 6'd45 - sum;
       b[32:1]<=a[32:1]; end
       default:  begin b[36:1]<=a[36:1]; end
    
  endcase
  end
endmodule
 ///module fullhouse///
module fullhouse( a_out,a,clk,rst,start);
  input [81*4:1] a;
    output reg [81*4:1] a_out;
    reg [81*4:1] b;
  reg [81*4:1] colmat;
  wire rept;
  parameter s0=3'd0,s1=3'd1,s2=3'd2,s3=3'd3,s4=3'd4,s5=3'd5,s6=3'd6,s7=3'd7;
  reg [3:0] state, nstate;
  reg assigning;
  input clk, rst,start;
  reg [36:1] fi1;
  reg [36:1] fo1;
  reg [36:1] fi2;
  reg [36:1] fo2;
  reg [36:1] fi3;
  reg [36:1] fo3;
  reg [36:1] fi4;
  reg [36:1] fo4;
  reg [36:1] fi5;
  reg [36:1] fo5;
  reg [36:1] fi6;
  reg [36:1] fo6;
  reg [36:1] fi7;
  reg [36:1] fo7;
  reg [36:1] fi8;
  reg [36:1] fo8;
  reg [36:1] fi9;
  reg [36:1] fo9;
  reg detection;
  reg [324:1] in;
  spacechk modl ( detection, in);
  
  
  reg fullrow, fullcol, fullbox, loadreg, asinput,resetf;
  genvar i,j;
  
  
  
    always @(posedge clk, negedge rst) begin
    if (~rst) 
      state<=s0;
  else 
    state<=nstate;
  end
 

  always @(state)
    begin
      case(state)
        s0: begin nstate=s1 ;loadreg=1; end
        
      s1: begin
           
            nstate<=s2;
            fi1<=b[36:1];
            fi2<=b[72:37];
            fi3<=b[108:73];
            fi4<=b[144:109];
            fi5<=b[180:145];
            fi6<=b[216:181];
            fi7<=b[252:217];
            fi8<=b[288:253];
            fi9<=b[324:289];
            fullrow=1'b1;
            
            end
        s2:begin
             nstate<=s3;
          fi1<={b[292:289],b[256:253],b[220:217],b[184:181],b[148:145],b[112:109],b[76:73],b[40:37],b[4:1]};
          fi2<={b[296:293],b[260:257],b[224:221],b[188:185],b[152:149],b[116:113],b[80:77],b[44:41],b[8:5]};
          fi3<={b[300:297],b[264:261],b[228:225],b[192:189],b[156:153],b[120:117],b[84:81],b[48:45],b[12:9]};
          fi4<={b[304:301],b[268:265],b[232:229],b[196:193],b[160:157],b[124:121],b[88:85],b[52:49],b[16:13]};
          fi5<={b[308:305],b[272:269],b[236:233],b[200:197],b[164:161],b[128:125],b[92:89],b[56:53],b[20:17]};
          fi6<={b[312:309],b[276:273],b[240:237],b[204:201],b[168:165],b[132:129],b[96:93],b[60:57],b[24:21]};
          fi7<={b[316:313],b[280:277],b[244:241],b[208:205],b[172:169],b[136:133],b[100:97],b[64:61],b[28:25]};
          fi8<={b[320:317],b[284:281],b[248:245],b[212:209],b[176:173],b[140:137],b[104:101],b[68:65],b[32:29]};
          fi9<={b[324:321],b[288:285],b[252:249],b[216:213],b[180:177],b[144:141],b[108:105],b[72:69],b[36:33]};
             fullcol=1'b1;
             end
          
        s3:begin
             nstate<=s4;
          fi1<={b[84:73],b[48:37],b[12:1]};
          fi2<={b[96:85],b[60:49],b[24:13]};
          fi3<={b[108:97],b[72:61],b[36:25]};
          fi4<={b[192:181],b[156:145],b[120:109]};
          fi5<={b[204:193],b[168:157],b[132:121]};
          fi6<={b[216:205],b[180:169],b[144:133]};
          fi7<={b[300:289],b[264:253],b[228:217]};
          fi8<={b[312:301],b[276:265],b[240:229]};
          fi9<={b[324:313],b[288:277],b[252:241]};
             fullbox=1;
             end
        
        s4: begin
            nstate<=s5;
            asinput=1'b1;
            end
        s5:begin
              
          if(detection) begin  nstate<=s1; end
          else nstate<=s6;
        end
         
        s6: assigning=1'b1;
     
        
      endcase
    end
  
  filler M1(fo1,fi1);
  filler M2(fo2,fi2);
  filler M3(fo3,fi3);
  filler M4(fo4,fi4);
  filler M5(fo5,fi5);
  filler M6(fo6,fi6);
  filler M7(fo7,fi7);
  filler M8(fo8,fi8);
  filler M9(fo9,fi9);
  always@(posedge clk)
    begin
          
      if (loadreg )
        begin
          
          b[324:1]<=a[324:1];
          loadreg=1'b0;
        end
      if (fullrow)
        begin
          
          b[36:1]<=fo1 ;
          b[72:37]<=fo2 ;
          b[108:73]<=fo3 ;
          b[144:109]<=fo4 ;
          b[180:145]<=fo5 ;
          b[216:181]<=fo6 ;
          b[252:217]<=fo7 ;
          b[288:253]<=fo8 ;
          b[324:289]<=fo9 ;
          fullrow=1'b0;
        end
      if (fullcol)
       begin
         {b[292:289],b[256:253],b[220:217],b[184:181],b[148:145],b[112:109],b[76:73],b[40:37],b[4:1]}<=fo1  ;
         {b[296:293],b[260:257],b[224:221],b[188:185],b[152:149],b[116:113],b[80:77],b[44:41],b[8:5]}<=fo2  ;
         {b[300:297],b[264:261],b[228:225],b[192:189],b[156:153],b[120:117],b[84:81],b[48:45],b[12:9]}<=fo3 ;
         {b[304:301],b[268:265],b[232:229],b[196:193],b[160:157],b[124:121],b[88:85],b[52:49],b[16:13]}<=fo4;
         {b[308:305],b[272:269],b[236:233],b[200:197],b[164:161],b[128:125],b[92:89],b[56:53],b[20:17]}<=fo5;
         {b[312:309],b[276:273],b[240:237],b[204:201],b[168:165],b[132:129],b[96:93],b[60:57],b[24:21]}<=fo6;
         {b[316:313],b[280:277],b[244:241],b[208:205],b[172:169],b[136:133],b[100:97],b[64:61],b[28:25]}<=fo7 ;
         {b[320:317],b[284:281],b[248:245],b[212:209],b[176:173],b[140:137],b[104:101],b[68:65],b[32:29]}<=fo8;
         {b[324:321],b[288:285],b[252:249],b[216:213],b[180:177],b[144:141],b[108:105],b[72:69],b[36:33]}<=fo9;
         fullcol=1'b0;
       end
      if(fullbox)
        begin
          {b[84:73],b[48:37],b[12:1]}<=fo1;
          {b[96:85],b[60:49],b[24:13]}<=fo2;
          {b[108:97],b[72:61],b[36:25]}<=fo3;
          {b[192:181],b[156:145],b[120:109]}<=fo4;
          {b[204:193],b[168:157],b[132:121]}<=fo5;
          {b[216:205],b[180:169],b[144:133]}<=fo6;
          {b[300:289],b[264:253],b[228:217]}<=fo7;
          {b[312:301],b[276:265],b[240:229]}<=fo8;
          {b[324:313],b[288:277],b[252:241]}<=fo9;
          fullbox=1'b0;
          
        end
      if(asinput)begin 
        in<=b;
        asinput=1'b0;
       
       end
      
      if (assigning)
        begin
          assign a_out=b;
        end
    end
              
endmodule


// Code your design here
// Code your design here
// Code your design here
module spacechk ( val, a);
  input  [324:1] a;
  output val;
  genvar i,j;
  reg [9:1] countr;
  reg [9:1]  countc,countb;
  wire [3:0] b,c,d,e,f,g,h,k,l,m,n,o,p,q,r,s,t,u,v,w,x,y,z,pp,sy,wr,rr;
  wire [4:1] trail= a[324:321] ;
  
  assign  b= !a[36:33]+ !a[32:29]+ !a[28:25] + !a[24:21] + !a[20:17] + !a[16:13] + !a[12:9] +!a[8:5] +!a[4:1];
  assign  c= !a[72:69]+ !a[68:65]+ !a[64:61] + !a[60:57] + !a[56:53] + !a[52:49] + !a[48:45]+!a[44:41] +!a[40:37];
  assign  d= !a[108:105]+ !a[104:101] + !a[100:97]  + !a[96:93]   + !a[92:89]  + !a[88:85]  + !a[84:81]   + !a[80:77]   + !a[76:73];
  assign  e= !a[144:141]+ !a[140:137] + !a[136:133] + !a[132:129] + !a[128:125]+ !a[124:121]+  !a[120:117]+ !a[116:113] + !a[112:109];
  assign  f= !a[180:177]+ !a[176:173] + !a[172:169] + !a[168:165] + !a[164:161]+ !a[160:157]+  !a[156:153]+ !a[152:149] + !a[148:145];
  assign  g= !a[216:213]+ !a[212:209] + !a[208:205] + !a[204:201] + !a[200:197]+ !a[196:193]+  !a[192:189]+ !a[188:185] + !a[184:181];
  assign  h= !a[252:249]+ !a[248:245] + !a[244:241] + !a[240:237] + !a[236:233]+ !a[232:229]+  !a[228:225]+ !a[224:221] + !a[220:217];
  assign  k= !a[288:285]+ !a[284:281] + !a[280:277] + !a[276:273] + !a[272:269]+ !a[268:265]+  !a[264:261]+ !a[260:257] + !a[256:253];
  assign  l= !a[324:321]+ !a[320:317] + !a[316:313] + !a[312:309] + !a[308:305]+ !a[304:301]+  !a[300:297]+ !a[296:293] + !a[292:289];
  
  assign  m= !a[292:289] + !a[256:253]+ !a[220:217]+ !a[184:181]+ !a[148:145]+ !a[112:109]+ !a[76:73]   + !a[40:37]+ !a[4:1];
  assign  n= !a[296:293] + !a[260:257]+ !a[224:221]+ !a[188:185]+ !a[152:149]+ !a[116:113]+ !a[80:77]   + !a[44:41]+ !a[8:5];
  assign  o= !a[300:297] + !a[264:261]+ !a[228:225]+ !a[192:189]+ !a[156:153]+ !a[120:117]+ !a[84:81]   + !a[48:45]+ !a[12:9];
  assign  p= !a[304:301] + !a[268:265]+ !a[232:229]+ !a[196:193]+ !a[160:157]+ !a[124:121]+ !a[88:85]   + !a[52:49]+ !a[16:13];
  assign  q= !a[308:305] + !a[272:269]+ !a[236:233]+ !a[200:197]+ !a[164:161]+ !a[128:125]+ !a[92:89]   + !a[56:53]+ !a[20:17];       
  assign  r= !a[312:309] + !a[276:273]+ !a[240:237]+ !a[204:201]+ !a[168:165]+ !a[132:129]+ !a[96:93]   + !a[60:57]+ !a[24:21];
  assign  s= !a[316:313] + !a[280:277]+ !a[244:241]+ !a[208:205]+ !a[172:169]+ !a[136:133]+ !a[100:97]  + !a[64:61]+ !a[28:25];
  assign  t= !a[320:317] + !a[284:281]+ !a[248:245]+ !a[212:209]+ !a[176:173]+ !a[140:137]+ !a[104:101] + !a[68:65]+ !a[32:29];
  assign  u= !a[324:321] + !a[288:285]+ !a[252:249]+ !a[216:213]+ !a[180:177]+ !a[144:141]+ !a[108:105] + !a[72:69]+ !a[36:33];
   
  assign  v=  !a[84:81]  + !a[80:77]  + !a[76:73]  + !a[40:37]  + !a[44:41]  + !a[48:45]  + !a[12:9]   + !a[8:5]    + !a[4:1];
  assign  w=  !a[96:93]  + !a[92:89]  + !a[88:85]  + !a[60:57]  + !a[56:53]  + !a[52:49]  + !a[24:21]  + !a[20:17]  + !a[16:13];
  assign  x=  !a[108:105]+ !a[104:101]+ !a[100:97] + !a[72:69]  + !a[68:65]  + !a[64:61]  + !a[36:33]  + !a[32:29]  + !a[28:25];
  assign  y=  !a[192:189]+ !a[188:185]+ !a[184:181]+ !a[156:153]+ !a[152:149]+ !a[148:145]+ !a[120:117]+ !a[116:113]+ !a[112:109];
  assign  z=  !a[132:129]+ !a[128:125]+ !a[124:121]+ !a[168:165]+ !a[164:161]+ !a[160:157]+ !a[204:201]+ !a[200:197]+ !a[196:193];
  assign  pp= !a[216:213]+ !a[212:209]+ !a[208:205]+ !a[180:177]+ !a[176:173]+ !a[172:169]+ !a[144:141]+ !a[140:137]+ !a[136:133];
  assign  sy= !a[300:297]+ !a[296:293]+ !a[292:289]+ !a[264:261]+ !a[260:257]+ !a[256:253]+ !a[228:225]+ !a[224:221]+ !a[220:217];
  assign  wr= !a[312:309]+ !a[308:305]+ !a[304:301]+ !a[276:273]+ !a[272:269]+ !a[268:265]+ !a[240:237]+ !a[236:233]+ !a[232:229];
  assign  rr= !a[324:321]+ !a[320:317]+ !a[316:313]+ !a[252:249]+ !a[248:245]+ !a[244:241]+ !a[238:235]+ !a[234:231]+ !a[230:227];
         
  
  assign val=  (b==1)| (c==1)| (d==1)| (e==1)| (f==1)| (g==1)| (h==1)| (k==1)| (l==1)| (m==1)| (n==1)| (o==1)| (p==1)| (q==1)| (r==1)| (s==1)| (t==1)| (u==1)| (v==1)| (x==1) | (y==1)| (z==1)| (wr==1)| (pp==1)| (rr==1)| (s==1)| (w==1);
endmodule



